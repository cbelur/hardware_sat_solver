`timescale 1ns / 1ps 
import common::*;
module top_test();
logic clock, reset, load;
logic[number_literal-1:0] i;
logic ended, sat;
logic[number_literal-1:0] model;
top test1(clock, reset, load, i, ended, sat, model);
always
begin
clock=1'b1; #50; clock=1'b0; #50;
end
initial
begin
reset=1'b1; load <= 1'b0;
#60;
reset=1'b0; load <= 1'b1;)





i <= 30'b110000000000000000000000000000; #100; 
i <= 30'b000000000000000000000000000000; #100; 
i <= 30'b101000000000000000000000000000; #100; 
i <= 30'b000000000000000000000000000000; #100; 
i <= 30'b010000000000000000000000000000; #100; 
i <= 30'b101000000000000000000000000000; #100; 
i <= 30'b000000000000000000000000000000; #100; 
i <= 30'b011000000000000000000000000000; #100; 
i <= 30'b011000000000000000000000000000; #100; 
i <= 30'b100000000000000000000000000000; #100; 
i <= 30'b100000000000000000000000000000; #100; 
i <= 30'b000100000000000000000000000000; #100; 
i <= 30'b010000000000000000000000000000; #100; 
i <= 30'b000100000000000000000000000000; #100; 
i <= 30'b000100000000000000000000000000; #100; 
i <= 30'b110000000000000000000000000000; #100; 
i <= 30'b000000100000000000000000000000; #100; 
i <= 30'b000000000100000000000000000000; #100; 
i <= 30'b000000010000000000000000000000; #100; 
i <= 30'b000000000100000000000000000000; #100; 
i <= 30'b000000000100000000000000000000; #100; 
i <= 30'b000000110000000000000000000000; #100; 
i <= 30'b000000000000100000000000000000; #100; 
i <= 30'b000000000000000100000000000000; #100; 
i <= 30'b000000000000010000000000000000; #100; 
i <= 30'b000000000000000100000000000000; #100; 
i <= 30'b000000000000000100000000000000; #100; 
i <= 30'b000000000000110000000000000000; #100; 
i <= 30'b000000000000000000100000000000; #100; 
i <= 30'b000000000000000000000100000000; #100; 
i <= 30'b000000000000000000010000000000; #100; 
i <= 30'b000000000000000000000100000000; #100; 
i <= 30'b000000000000000000000100000000; #100; 
i <= 30'b000000000000000000110000000000; #100; 
i <= 30'b000000000000000000000000100000; #100; 
i <= 30'b000000000000000000000000000100; #100; 
i <= 30'b000000000000000000000000010000; #100; 
i <= 30'b000000000000000000000000000100; #100; 
i <= 30'b000000000000000000000000000100; #100; 
i <= 30'b000000000000000000000000110000; #100; 
i <= 30'b000000000000000000000000000000; #100; 
i <= 30'b000110000000000000000000000000; #100; 
i <= 30'b000110000000000000000000000000; #100; 
i <= 30'b000000000000000000000000000000; #100; 
i <= 30'b000000000000000000000000000000; #100; 
i <= 30'b000000000110000000000000000000; #100; 
i <= 30'b000000000110000000000000000000; #100; 
i <= 30'b000000000000000000000000000000; #100; 
i <= 30'b000000000000000000000000000000; #100; 
i <= 30'b000000000000000110000000000000; #100; 
i <= 30'b000000000000000110000000000000; #100; 
i <= 30'b000000000000000000000000000000; #100; 
i <= 30'b000000000000000000000000000000; #100; 
i <= 30'b000000000000000000000110000000; #100; 
i <= 30'b000000000000000000000110000000; #100; 
i <= 30'b000000000000000000000000000000; #100; 
i <= 30'b000000000000000000000000000000; #100; 
i <= 30'b000000000000000000000000000110; #100; 
i <= 30'b000000000000000000000000000110; #100; 
i <= 30'b000000000000000000000000000000; #100; 
i <= 30'b000000000000000000000000000000; #100; 
i <= 30'b001001000000000000000000000000; #100; 
i <= 30'b001001000000000000000000000000; #100; 
i <= 30'b000000000000000000000000000000; #100; 
i <= 30'b000000000000000000000000000000; #100; 
i <= 30'b000000001001000000000000000000; #100; 
i <= 30'b000000001001000000000000000000; #100; 
i <= 30'b000000000000000000000000000000; #100; 
i <= 30'b000000000000000000000000000000; #100; 
i <= 30'b000000000000001001000000000000; #100; 
i <= 30'b000000000000001001000000000000; #100; 
i <= 30'b000000000000000000000000000000; #100; 
i <= 30'b000000000000000000000000000000; #100; 
i <= 30'b000000000000000000001001000000; #100; 
i <= 30'b000000000000000000001001000000; #100; 
i <= 30'b000000000000000000000000000000; #100; 
i <= 30'b000000000000000000000000000000; #100; 
i <= 30'b000000000000000000000000001001; #100; 
i <= 30'b000000000000000000000000001001; #100; 
i <= 30'b000000000000000000000000000000; #100; 
i <= 30'b000000010000000000000000000000; #100; 
i <= 30'b000010000000000000000000000000; #100; 
i <= 30'b000010000000000000000000000000; #100; 
i <= 30'b000000010000000000000000000000; #100; 
i <= 30'b000000001000000000000000000000; #100; 
i <= 30'b000001000000000000000000000000; #100; 
i <= 30'b000001000000000000000000000000; #100; 
i <= 30'b000000001000000000000000000000; #100; 
i <= 30'b000000000000010000000000000000; #100; 
i <= 30'b000000000010000000000000000000; #100; 
i <= 30'b000000000010000000000000000000; #100; 
i <= 30'b000000000000010000000000000000; #100; 
i <= 30'b000000000000001000000000000000; #100; 
i <= 30'b000000000001000000000000000000; #100; 
i <= 30'b000000000001000000000000000000; #100; 
i <= 30'b000000000000001000000000000000; #100; 
i <= 30'b000000000000000000010000000000; #100; 
i <= 30'b000000000000000010000000000000; #100; 
i <= 30'b000000000000000010000000000000; #100; 
i <= 30'b000000000000000000010000000000; #100; 
i <= 30'b000000000000000000001000000000; #100; 
i <= 30'b000000000000000001000000000000; #100; 
i <= 30'b000000000000000001000000000000; #100; 
i <= 30'b000000000000000000001000000000; #100; 
i <= 30'b000000000000000000000000010000; #100; 
i <= 30'b000000000000000000000010000000; #100; 
i <= 30'b000000000000000000000010000000; #100; 
i <= 30'b000000000000000000000000010000; #100; 
i <= 30'b000000000000000000000000001000; #100; 
i <= 30'b000000000000000000000001000000; #100; 
i <= 30'b000000000000000000000001000000; #100; 
i <= 30'b000000000000000000000000001000; #100; 
i <= 30'b000000000000000000000000000000; #100; 
i <= 30'b010000000000000000000000000000; #100; 
i <= 30'b000000000000000000000000000000; #100; 
i <= 30'b001000000000000000000000000000; #100; 
i <= 30'b000000000000000000000000000010; #100; 
i <= 30'b000000000000000000000000000000; #100; 
i <= 30'b000000000000000000000000000001; #100; 
i <= 30'b000000000000000000000000000000; #100; 
load <= 1'b0; 
end
endmodule
